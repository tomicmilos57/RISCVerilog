module instruction_register(clk, in, valid, state, out, instruction);

// ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==
//  Ports
// ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==

input        clk;
input [31:0] in;
input        valid;
input        state;
input [31:0] out;
input [31:0] instruction;

// ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==
//  Combinational Logic
// ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==

reg [31:0] r_IR;
assign out = r_IR;

reg[31:0] r_instruction;
assign instruction = r_instruction;

wire FETCH = state == 1'h0;
wire EXECUTE = state == 1'h1;

// ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==
//  Sequential Logic
// ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==  ==

always @(posedge clk) begin
  if(FETCH & valid) begin
    r_IR <= in;
    case (in)
      // R-type instructions (opcode = 0110011)
      32'b0000000_?????_?????_000_?????_0110011: r_instruction = 32'd0;  // ADD
      32'b0100000_?????_?????_000_?????_0110011: r_instruction = 32'd1;  // SUB
      32'b0000000_?????_?????_001_?????_0110011: r_instruction = 32'd2;  // SLL
      32'b0000000_?????_?????_010_?????_0110011: r_instruction = 32'd3;  // SLT
      32'b0000000_?????_?????_011_?????_0110011: r_instruction = 32'd4;  // SLTU
      32'b0000000_?????_?????_100_?????_0110011: r_instruction = 32'd5;  // XOR
      32'b0000000_?????_?????_101_?????_0110011: r_instruction = 32'd6;  // SRL
      32'b0100000_?????_?????_101_?????_0110011: r_instruction = 32'd7;  // SRA
      32'b0000000_?????_?????_110_?????_0110011: r_instruction = 32'd8;  // OR
      32'b0000000_?????_?????_111_?????_0110011: r_instruction = 32'd9;  // AND

      // Multiplication and Division instructions (RV32M, opcode = 0110011)
      32'b0000001_?????_?????_000_?????_0110011: r_instruction = 32'd10; // MUL
      32'b0000001_?????_?????_001_?????_0110011: r_instruction = 32'd11; // MULH
      32'b0000001_?????_?????_010_?????_0110011: r_instruction = 32'd12; // MULHSU
      32'b0000001_?????_?????_011_?????_0110011: r_instruction = 32'd13; // MULHU
      32'b0000001_?????_?????_100_?????_0110011: r_instruction = 32'd14; // DIV
      32'b0000001_?????_?????_101_?????_0110011: r_instruction = 32'd15; // DIVU
      32'b0000001_?????_?????_110_?????_0110011: r_instruction = 32'd16; // REM
      32'b0000001_?????_?????_111_?????_0110011: r_instruction = 32'd17; // REMU

      // I-type instructions (opcode = 0010011)
      32'b????????????_?????_000_?????_0010011: r_instruction = 32'd18; // ADDI
      32'b????????????_?????_010_?????_0010011: r_instruction = 32'd19; // SLTI
      32'b????????????_?????_011_?????_0010011: r_instruction = 32'd20; // SLTIU
      32'b????????????_?????_100_?????_0010011: r_instruction = 32'd21; // XORI
      32'b????????????_?????_110_?????_0010011: r_instruction = 32'd22; // ORI
      32'b????????????_?????_111_?????_0010011: r_instruction = 32'd23; // ANDI
      32'b0000000_?????_?????_001_?????_0010011: r_instruction = 32'd24; // SLLI
      32'b0000000_?????_?????_101_?????_0010011: r_instruction = 32'd25; // SRLI
      32'b0100000_?????_?????_101_?????_0010011: r_instruction = 32'd26; // SRAI

      // Load instructions (opcode = 0000011)
      32'b????????????_?????_000_?????_0000011: r_instruction = 32'd27; // LB
      32'b????????????_?????_001_?????_0000011: r_instruction = 32'd28; // LH
      32'b????????????_?????_010_?????_0000011: r_instruction = 32'd29; // LW
      32'b????????????_?????_100_?????_0000011: r_instruction = 32'd30; // LBU
      32'b????????????_?????_101_?????_0000011: r_instruction = 32'd31; // LHU

      // S-type instructions (opcode = 0100011)
      32'b????????????_?????_000_?????_0100011: r_instruction = 32'd32; // SB
      32'b????????????_?????_001_?????_0100011: r_instruction = 32'd33; // SH
      32'b????????????_?????_010_?????_0100011: r_instruction = 32'd34; // SW

      // B-type instructions (opcode = 1100011)
      32'b????????????_?????_000_?????_1100011: r_instruction = 32'd35; // BEQ
      32'b????????????_?????_001_?????_1100011: r_instruction = 32'd36; // BNE
      32'b????????????_?????_100_?????_1100011: r_instruction = 32'd37; // BLT
      32'b????????????_?????_101_?????_1100011: r_instruction = 32'd38; // BGE
      32'b????????????_?????_110_?????_1100011: r_instruction = 32'd39; // BLTU
      32'b????????????_?????_111_?????_1100011: r_instruction = 32'd40; // BGEU

      // J-type instructions (opcode = 1101111)
      32'b????????????????????_?????_1101111: r_instruction = 32'd41; // JAL

      // I-type instructions (opcode = 1100111)
      32'b????????????_?????_000_?????_1100111: r_instruction = 32'd42; // JALR

      // U-type instructions (opcode = 0110111)
      32'b????????????????????_?????_0110111: r_instruction = 32'd43; // LUI

      // U-type instructions (opcode = 0010111)
      32'b????????????????????_?????_0010111: r_instruction = 32'd44; // AUIPC

      default: r_instruction = 32'd45; // Unknown or unsupported instruction
    endcase
    //Clear r_IR if EXECUTE state ?
  end
end

endmodule

